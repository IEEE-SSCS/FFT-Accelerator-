module cordic #(
parameter data_width=8
)
(
input logic clk,nrst,
input  logic [data_width-1:0] in_real,in_img,
input  logic [data_width-1:0] FA_sgn,
output logic [data_width-1:0] out_real,out_img
);










endmodule